module XTEA_DEC (
    ports
);
    
endmodule